Changes made in repo2
